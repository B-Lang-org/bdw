
module Empty(CLK, RST);
   input     CLK;
   input     RST;


endmodule

